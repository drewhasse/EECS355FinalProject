library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity tank_game is
  port (
  );
end entity;

architecture structural of tank_game is

begin

end architecture;
